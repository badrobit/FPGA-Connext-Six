module game_board();

// 19x19 array of 4 bit registers. 
// reg = X | XXX 
reg [3:0] game_board [0:18] [0:18];

endmodule