module controller
(
	input 		clock_50, 
	input [3:0]	Key,

	//output - to serial :) 
);

endmodule 