module controller();



endmodule 